// *********************************************************
// Program: hours.sv
// Description: counts hours on the clock
// Author: Jeffrey Noe
// Due: 6/8/2018
// *********************************************************

module hours (
      input                   clkMSec,
      input                   resetN,
      input                   milTime,
      output logic            amPm,
      output logic [4:0]      hour
      );


endmodule
