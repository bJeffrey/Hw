// *********************************************************
// Program: minutes.sv
// Description: counts minutes on the clock
// Author: Jeffrey Noe
// Due: 6/8/2018
// *********************************************************

module minutes (
      input                   clkMSec,
      input                   resetN,
      output logic            changeHour,
      output logic [5:0]      min
      );


endmodule
